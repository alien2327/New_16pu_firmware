interface dc1884a_int;
    logic [ 1:0] data_clk_in_p;
    logic [ 1:0] data_clk_in_n;
    logic [ 1:0] frame_in_p;
    logic [ 1:0] frame_in_n;
    logic [15:0] data_in_p;
    logic [15:0] data_in_n;
endinterface

module 16pu_main #(
    parameter dummy = 0
) (

);



endmodule