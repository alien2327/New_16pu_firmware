module sitcp_wrap(

);

endmodule