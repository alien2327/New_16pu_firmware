module 16pu_main #(
    parameter dummy = 0
) (

);



endmodule