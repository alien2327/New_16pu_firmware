module deepfifo_wrap(

);

endmodule