module lcd_wrap(

);

endmodule