interface rbcp_int;
    logic        RBCP_WE;
    logic        RBCP_RE;
    logic [ 7:0] RBCP_WD;
    logic [31:0] RBCP_ADDR;
    logic [ 7:0] RBCP_RD;
    logic		 RBCP_ACK;
endinterface

module sitcp_wrap(

);

endmodule