module adc_capture_wrap(

);

endmodule